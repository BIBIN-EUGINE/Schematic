-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Friday, May 24, 2019 11:25:38 Eastern Daylight Time

